CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 80 1364 699
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 46 632 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9672 0 0
2
45910.9 0
0
13 Logic Switch~
5 52 527 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7876 0 0
2
45910.9 0
0
13 Logic Switch~
5 176 421 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6369 0 0
2
45910.9 0
0
13 Logic Switch~
5 178 297 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9172 0 0
2
45910.9 0
0
13 Logic Switch~
5 180 276 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
45910.9 0
0
13 Logic Switch~
5 214 177 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3820 0 0
2
45910.9 0
0
13 Logic Switch~
5 208 95 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7678 0 0
2
45910.9 0
0
14 Logic Display~
6 496 564 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
961 0 0
2
45910.9 0
0
9 2-In NOR~
219 348 576 0 3 22
0 4 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3178 0 0
2
45910.9 0
0
9 2-In NOR~
219 213 617 0 3 22
0 7 5 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3409 0 0
2
45910.9 0
0
9 2-In NOR~
219 214 543 0 3 22
0 6 7 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3951 0 0
2
45910.9 0
0
9 2-In NOR~
219 112 579 0 3 22
0 6 5 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8885 0 0
2
45910.9 0
0
14 Logic Display~
6 399 417 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3780 0 0
2
45910.9 0
0
9 2-In NOR~
219 263 422 0 3 22
0 8 8 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9265 0 0
2
45910.9 0
0
14 Logic Display~
6 451 276 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9442 0 0
2
45910.9 0
0
9 2-In NOR~
219 375 288 0 3 22
0 13 13 10
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9424 0 0
2
45910.9 0
0
9 2-In NOR~
219 224 286 0 3 22
0 12 11 13
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9968 0 0
2
45910.9 0
0
9 2-In NOR~
219 414 127 0 3 22
0 18 17 14
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9281 0 0
2
45910.9 0
0
9 2-In NOR~
219 277 176 0 3 22
0 15 15 17
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8464 0 0
2
45910.9 0
0
9 2-In NOR~
219 277 96 0 3 22
0 16 16 18
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7168 0 0
2
45910.9 0
0
14 Logic Display~
6 476 105 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3171 0 0
2
45910.9 0
0
24
3 1 2 0 0 4224 0 9 8 0 0 5
387 576
484 576
484 590
496 590
496 582
2 3 3 0 0 4224 0 9 10 0 0 4
335 585
260 585
260 617
252 617
3 1 4 0 0 4224 0 11 9 0 0 4
253 543
327 543
327 567
335 567
2 1 5 0 0 4224 0 10 1 0 0 4
200 626
72 626
72 632
58 632
1 1 6 0 0 4224 0 11 2 0 0 4
201 534
78 534
78 527
64 527
2 1 5 0 0 0 0 12 1 0 0 4
99 588
67 588
67 632
58 632
1 1 6 0 0 0 0 12 2 0 0 4
99 570
73 570
73 527
64 527
3 0 7 0 0 4096 0 12 0 0 9 2
151 579
192 579
2 1 7 0 0 8320 0 11 10 0 0 4
201 552
192 552
192 608
200 608
1 0 8 0 0 4224 0 3 0 0 12 4
188 421
237 421
237 422
242 422
3 1 9 0 0 4224 0 14 13 0 0 5
302 422
387 422
387 443
399 443
399 435
1 2 8 0 0 0 0 14 14 0 0 4
250 413
242 413
242 431
250 431
3 1 10 0 0 4224 0 16 15 0 0 5
414 288
439 288
439 302
451 302
451 294
1 2 11 0 0 4224 0 4 17 0 0 4
190 297
203 297
203 295
211 295
1 1 12 0 0 4224 0 5 17 0 0 4
192 276
203 276
203 277
211 277
3 0 13 0 0 4224 0 17 0 0 17 2
263 286
354 286
1 2 13 0 0 0 0 16 16 0 0 4
362 279
354 279
354 297
362 297
3 1 14 0 0 4240 0 18 21 0 0 3
453 127
476 127
476 123
1 0 15 0 0 4224 0 6 0 0 23 2
226 177
255 177
1 0 16 0 0 4224 0 7 0 0 24 2
220 95
255 95
3 2 17 0 0 4224 0 19 18 0 0 5
316 176
392 176
392 141
401 141
401 136
3 1 18 0 0 8320 0 20 18 0 0 6
316 96
316 97
392 97
392 116
401 116
401 118
1 2 15 0 0 0 0 19 19 0 0 4
264 167
255 167
255 185
264 185
1 2 16 0 0 0 0 20 20 0 0 6
264 87
256 87
256 88
255 88
255 105
264 105
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
176 476 355 500
181 480 349 496
21 NOR GATE AS XNOR GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
230 351 361 375
235 355 355 371
15 NOR gate as NOT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
264 220 427 244
269 224 421 240
19 NOR Gate as OR Gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
249 25 420 49
254 29 414 45
20 NOR Gate as AND Gate
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
