CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 30 70 10
337 149 1168 551
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
505 245 618 342
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 46 859 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9672 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 43 715 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 101 548 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6369 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 103 409 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 95 329 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7100 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 71 222 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3820 0 0
2
5.90184e-315 0
0
13 Logic Switch~
5 73 153 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7678 0 0
2
5.90184e-315 0
0
14 Logic Display~
6 517 739 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 414 766 0 3 22
0 4 3 2
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3178 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 250 846 0 3 22
0 5 6 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3409 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 248 723 0 3 22
0 7 5 4
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3951 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 151 777 0 3 22
0 7 6 5
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
8885 0 0
2
5.90184e-315 0
0
14 Logic Display~
6 460 541 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 284 548 0 3 22
0 9 9 8
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9265 0 0
2
5.90184e-315 0
0
14 Logic Display~
6 557 354 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 374 363 0 3 22
0 11 12 10
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9424 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 253 413 0 3 22
0 13 13 12
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
9968 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 251 341 0 3 22
0 14 14 11
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
9281 0 0
2
5.90184e-315 0
0
14 Logic Display~
6 430 163 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 330 180 0 3 22
0 16 16 15
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7168 0 0
2
5.90184e-315 0
0
10 2-In NAND~
219 183 180 0 3 22
0 18 17 16
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3171 0 0
2
5.90184e-315 0
0
24
3 1 2 0 0 4224 0 9 8 0 0 3
441 766
517 766
517 757
3 2 3 0 0 4224 0 10 9 0 0 4
277 846
385 846
385 775
390 775
3 1 4 0 0 4224 0 11 9 0 0 4
275 723
384 723
384 757
390 757
0 2 5 0 0 4096 0 0 11 5 0 3
219 777
219 732
224 732
3 1 5 0 0 8320 0 12 10 0 0 4
178 777
220 777
220 837
226 837
1 2 6 0 0 4240 0 1 10 0 0 3
58 859
226 859
226 855
1 1 7 0 0 8320 0 2 11 0 0 3
55 715
55 714
224 714
2 1 6 0 0 0 0 12 1 0 0 3
127 786
58 786
58 859
1 1 7 0 0 0 0 2 12 0 0 3
55 715
55 768
127 768
3 1 8 0 0 4224 0 14 13 0 0 5
311 548
448 548
448 567
460 567
460 559
1 0 9 0 0 4224 0 3 0 0 12 4
113 548
247 548
247 549
252 549
1 2 9 0 0 0 0 14 14 0 0 4
260 539
252 539
252 557
260 557
3 1 10 0 0 4224 0 16 15 0 0 5
401 363
545 363
545 380
557 380
557 372
3 1 11 0 0 4224 0 18 16 0 0 4
278 341
342 341
342 354
350 354
3 2 12 0 0 4224 0 17 16 0 0 4
280 413
342 413
342 372
350 372
1 0 13 0 0 4224 0 4 0 0 17 2
115 409
221 409
1 2 13 0 0 0 0 17 17 0 0 4
229 404
221 404
221 422
229 422
1 0 14 0 0 4224 0 5 0 0 19 4
107 329
214 329
214 341
219 341
1 2 14 0 0 0 0 18 18 0 0 4
227 332
219 332
219 350
227 350
3 1 15 0 0 8320 0 20 19 0 0 3
357 180
357 181
430 181
0 3 16 0 0 4224 0 0 21 22 0 2
306 180
210 180
1 2 16 0 0 0 0 20 20 0 0 2
306 171
306 189
1 2 17 0 0 4224 0 6 21 0 0 4
83 222
144 222
144 189
159 189
1 1 18 0 0 4224 0 7 21 0 0 4
85 153
144 153
144 171
159 171
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
734 161 871 176
749 173 855 184
15 HAMMAD RIAZ 075
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
236 89 419 113
243 94 411 110
21 NAND GATE TO AND GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
269 273 444 297
276 279 436 295
20 NAND GATE TO OR GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
223 481 406 505
230 487 398 503
21 NAND GATE TO NOT GATE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
101 627 260 651
108 633 252 649
18 NAND to Ex-OR Gate
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
